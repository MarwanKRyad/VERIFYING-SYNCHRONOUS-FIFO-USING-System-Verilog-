package shared_pkg;
int error_count=0;
int correct_count=0;
bit finished_signal=0;
endpackage 
